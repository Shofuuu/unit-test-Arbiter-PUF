`ifndef defined
`define defined

parameter C_LENGTH = 64; // Length of the multiplexer challenge inputs

`endif // defined